package spi_test_pkg;

  import uvm_pkg::*;
  import apb_agent_pkg::*;
  import spi_agent_pkg::*;
  import spi_env_pkg::*;
  import spi_seq_pkg::*;

  `include "uvm_macros.svh"  
  `include "spi_test.svh"
  
endpackage: spi_test_pkg
  
  